# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__a41o_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.025000 1.450000 2.355000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 0.440000 1.815000 1.550000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.845000 0.440000 1.315000 1.550000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.455000 1.550000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.450000 2.925000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.639400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 0.350000 3.715000 0.770000 ;
        RECT 3.385000 0.770000 4.185000 0.940000 ;
        RECT 3.855000 1.820000 4.185000 2.980000 ;
        RECT 4.015000 0.940000 4.185000 1.820000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  1.720000 1.445000 1.890000 ;
      RECT 0.115000  1.890000 0.445000 2.980000 ;
      RECT 0.150000  0.085000 0.480000 1.010000 ;
      RECT 0.615000  2.060000 0.945000 3.245000 ;
      RECT 1.115000  1.890000 1.445000 1.950000 ;
      RECT 1.115000  1.950000 2.625000 2.120000 ;
      RECT 1.115000  2.120000 1.445000 2.980000 ;
      RECT 1.615000  2.290000 2.125000 3.245000 ;
      RECT 2.230000  0.350000 2.560000 1.110000 ;
      RECT 2.230000  1.110000 3.845000 1.280000 ;
      RECT 2.295000  2.120000 2.625000 2.980000 ;
      RECT 2.790000  0.085000 3.120000 0.940000 ;
      RECT 2.795000  1.950000 3.265000 2.120000 ;
      RECT 2.795000  2.120000 3.125000 2.980000 ;
      RECT 3.095000  1.280000 3.845000 1.550000 ;
      RECT 3.095000  1.550000 3.265000 1.950000 ;
      RECT 3.355000  2.270000 3.685000 3.245000 ;
      RECT 3.885000  0.085000 4.685000 0.600000 ;
      RECT 4.355000  1.820000 4.685000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__a41o_2
END LIBRARY
