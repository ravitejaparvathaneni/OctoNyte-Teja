# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__o211ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.685000 1.320000 4.695000 1.650000 ;
        RECT 4.365000 1.180000 4.695000 1.320000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 1.320000 3.445000 1.650000 ;
        RECT 2.435000 1.650000 3.235000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.350000 2.015000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 0.550000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.215200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.595000 0.890000 1.180000 ;
        RECT 0.595000 1.950000 3.285000 2.120000 ;
        RECT 0.595000 2.120000 0.925000 2.980000 ;
        RECT 0.720000 1.180000 0.890000 1.950000 ;
        RECT 1.495000 2.120000 1.825000 2.980000 ;
        RECT 2.955000 2.120000 3.285000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.130000  0.255000 2.330000 0.425000 ;
      RECT 0.130000  0.425000 0.380000 1.180000 ;
      RECT 0.145000  1.950000 0.395000 3.245000 ;
      RECT 1.060000  0.425000 2.330000 0.730000 ;
      RECT 1.060000  0.730000 1.390000 1.180000 ;
      RECT 1.125000  2.290000 1.295000 3.245000 ;
      RECT 1.560000  0.900000 1.890000 0.980000 ;
      RECT 1.560000  0.980000 4.160000 1.150000 ;
      RECT 1.560000  1.150000 1.890000 1.180000 ;
      RECT 2.025000  2.290000 2.275000 3.245000 ;
      RECT 2.505000  2.290000 2.755000 2.905000 ;
      RECT 2.505000  2.905000 3.655000 3.075000 ;
      RECT 2.560000  0.085000 2.890000 0.795000 ;
      RECT 3.070000  0.350000 3.240000 0.980000 ;
      RECT 3.420000  0.085000 3.750000 0.795000 ;
      RECT 3.485000  1.820000 4.685000 1.990000 ;
      RECT 3.485000  1.990000 3.655000 2.905000 ;
      RECT 3.855000  2.160000 4.185000 3.245000 ;
      RECT 3.935000  0.350000 4.160000 0.980000 ;
      RECT 4.330000  0.085000 4.685000 1.010000 ;
      RECT 4.355000  1.990000 4.685000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_hs__o211ai_2
END LIBRARY
