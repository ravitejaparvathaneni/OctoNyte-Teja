# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__dfstp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 0.980000 0.805000 1.990000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.119700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.680000 0.350000 11.010000 0.980000 ;
        RECT 10.680000 0.980000 12.835000 1.150000 ;
        RECT 11.175000 1.820000 12.835000 2.080000 ;
        RECT 11.175000 2.080000 11.455000 2.980000 ;
        RECT 12.015000 0.350000 12.345000 0.980000 ;
        RECT 12.125000 2.080000 12.835000 2.150000 ;
        RECT 12.125000 2.150000 12.355000 2.980000 ;
        RECT 12.605000 1.150000 12.835000 1.820000 ;
    END
  END Q
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  2.205000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.375000 1.550000 5.665000 1.595000 ;
        RECT 5.375000 1.595000 8.545000 1.735000 ;
        RECT 5.375000 1.735000 5.665000 1.780000 ;
        RECT 8.255000 1.550000 8.545000 1.595000 ;
        RECT 8.255000 1.735000 8.545000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.180000 1.775000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.115000  0.350000  0.365000 0.810000 ;
      RECT  0.115000  0.810000  0.285000 2.240000 ;
      RECT  0.115000  2.240000  1.795000 2.410000 ;
      RECT  0.115000  2.410000  0.365000 2.960000 ;
      RECT  0.545000  0.085000  0.795000 0.810000 ;
      RECT  0.565000  2.580000  0.895000 3.245000 ;
      RECT  0.975000  0.340000  1.435000 1.010000 ;
      RECT  0.975000  1.010000  1.145000 1.720000 ;
      RECT  0.975000  1.720000  2.275000 1.890000 ;
      RECT  0.975000  1.890000  1.455000 2.070000 ;
      RECT  1.575000  2.580000  1.905000 3.245000 ;
      RECT  1.615000  0.085000  1.865000 1.010000 ;
      RECT  1.625000  2.070000  2.615000 2.240000 ;
      RECT  1.945000  1.350000  2.275000 1.720000 ;
      RECT  2.045000  0.255000  3.115000 0.425000 ;
      RECT  2.045000  0.425000  2.215000 1.130000 ;
      RECT  2.105000  2.410000  2.275000 2.905000 ;
      RECT  2.105000  2.905000  3.795000 3.075000 ;
      RECT  2.445000  0.595000  2.775000 0.925000 ;
      RECT  2.445000  0.925000  2.615000 2.070000 ;
      RECT  2.445000  2.240000  2.615000 2.295000 ;
      RECT  2.445000  2.295000  2.945000 2.735000 ;
      RECT  2.785000  1.455000  3.115000 2.125000 ;
      RECT  2.945000  0.425000  3.115000 1.455000 ;
      RECT  3.115000  2.295000  3.455000 2.735000 ;
      RECT  3.285000  0.350000  3.535000 1.130000 ;
      RECT  3.285000  1.130000  4.135000 1.300000 ;
      RECT  3.285000  1.300000  3.455000 2.295000 ;
      RECT  3.625000  1.470000  3.795000 2.165000 ;
      RECT  3.625000  2.165000  4.685000 2.335000 ;
      RECT  3.625000  2.335000  3.795000 2.905000 ;
      RECT  3.965000  1.300000  4.135000 1.400000 ;
      RECT  3.965000  1.400000  5.025000 1.570000 ;
      RECT  3.985000  2.505000  4.345000 2.755000 ;
      RECT  3.985000  2.755000  4.155000 3.245000 ;
      RECT  4.025000  0.085000  4.420000 0.600000 ;
      RECT  4.115000  1.740000  5.025000 1.995000 ;
      RECT  4.305000  0.780000  5.050000 0.950000 ;
      RECT  4.305000  0.950000  4.590000 1.230000 ;
      RECT  4.515000  2.335000  4.685000 2.905000 ;
      RECT  4.515000  2.905000  5.510000 3.075000 ;
      RECT  4.590000  0.620000  5.050000 0.780000 ;
      RECT  4.770000  1.120000  5.025000 1.200000 ;
      RECT  4.770000  1.200000  6.135000 1.370000 ;
      RECT  4.770000  1.370000  5.025000 1.400000 ;
      RECT  4.855000  1.995000  5.025000 2.295000 ;
      RECT  4.855000  2.295000  5.170000 2.735000 ;
      RECT  5.195000  1.550000  5.635000 1.925000 ;
      RECT  5.340000  2.095000  6.475000 2.265000 ;
      RECT  5.340000  2.265000  5.510000 2.905000 ;
      RECT  5.670000  0.085000  6.000000 1.030000 ;
      RECT  5.680000  2.435000  5.940000 3.245000 ;
      RECT  5.805000  1.370000  6.135000 1.490000 ;
      RECT  6.305000  0.255000  7.375000 0.425000 ;
      RECT  6.305000  0.425000  6.475000 1.120000 ;
      RECT  6.305000  1.120000  6.695000 1.450000 ;
      RECT  6.305000  1.450000  6.475000 2.095000 ;
      RECT  6.590000  2.650000  7.265000 2.980000 ;
      RECT  6.645000  0.595000  7.035000 0.925000 ;
      RECT  6.670000  1.620000  7.035000 1.790000 ;
      RECT  6.670000  1.790000  6.840000 2.480000 ;
      RECT  6.670000  2.480000  7.715000 2.650000 ;
      RECT  6.865000  0.925000  7.035000 1.620000 ;
      RECT  7.045000  2.020000  7.375000 2.310000 ;
      RECT  7.205000  0.425000  7.375000 2.020000 ;
      RECT  7.545000  0.840000  9.450000 1.010000 ;
      RECT  7.545000  1.010000  7.875000 1.655000 ;
      RECT  7.545000  2.310000  9.110000 2.480000 ;
      RECT  7.885000  2.650000  8.055000 3.245000 ;
      RECT  7.935000  0.085000  8.950000 0.670000 ;
      RECT  8.185000  1.180000  8.515000 1.850000 ;
      RECT  8.255000  2.480000  8.585000 2.980000 ;
      RECT  8.780000  1.370000  9.110000 2.310000 ;
      RECT  8.780000  2.650000  9.030000 3.245000 ;
      RECT  9.120000  0.420000  9.450000 0.840000 ;
      RECT  9.230000  2.650000  9.560000 2.980000 ;
      RECT  9.280000  1.010000  9.450000 2.650000 ;
      RECT  9.680000  0.350000 10.010000 1.320000 ;
      RECT  9.680000  1.320000 11.995000 1.490000 ;
      RECT  9.755000  1.820000 10.005000 3.245000 ;
      RECT 10.180000  0.085000 10.510000 1.130000 ;
      RECT 10.205000  1.490000 11.995000 1.650000 ;
      RECT 10.205000  1.650000 10.535000 2.700000 ;
      RECT 10.725000  1.820000 11.005000 3.245000 ;
      RECT 11.180000  0.085000 11.845000 0.800000 ;
      RECT 11.625000  2.250000 11.955000 3.245000 ;
      RECT 12.515000  0.085000 12.845000 0.810000 ;
      RECT 12.525000  2.320000 12.855000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.580000  5.605000 1.750000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  1.580000  8.485000 1.750000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
  END
END sky130_fd_sc_hs__dfstp_4
END LIBRARY
