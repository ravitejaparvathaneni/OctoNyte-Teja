# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__dlygate4sd1_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.509700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.325000 0.355000 3.740000 1.120000 ;
        RECT 3.325000 1.815000 3.740000 3.060000 ;
        RECT 3.450000 1.120000 3.740000 1.815000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.095000  0.305000 0.410000 0.820000 ;
      RECT 0.095000  0.820000 1.305000 1.020000 ;
      RECT 0.095000  2.030000 1.305000 2.205000 ;
      RECT 0.095000  2.205000 0.400000 2.725000 ;
      RECT 0.575000  2.380000 0.905000 3.245000 ;
      RECT 0.585000  0.085000 0.915000 0.650000 ;
      RECT 0.975000  1.020000 1.305000 2.030000 ;
      RECT 1.415000  0.305000 1.720000 0.635000 ;
      RECT 1.415000  2.395000 1.720000 2.725000 ;
      RECT 1.475000  0.635000 1.720000 1.380000 ;
      RECT 1.475000  1.380000 2.740000 1.610000 ;
      RECT 1.475000  1.610000 1.720000 2.395000 ;
      RECT 1.985000  0.710000 2.345000 1.040000 ;
      RECT 1.985000  1.040000 3.155000 1.210000 ;
      RECT 1.985000  1.825000 3.155000 1.995000 ;
      RECT 1.985000  1.995000 2.345000 2.190000 ;
      RECT 2.825000  0.085000 3.155000 0.870000 ;
      RECT 2.825000  2.165000 3.155000 3.245000 ;
      RECT 2.910000  1.210000 3.155000 1.295000 ;
      RECT 2.910000  1.295000 3.280000 1.625000 ;
      RECT 2.910000  1.625000 3.155000 1.825000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_hs__dlygate4sd1_1
END LIBRARY
