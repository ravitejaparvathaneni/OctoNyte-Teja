# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__nand2b_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.363000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 1.115000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.780000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845000 1.300000 5.655000 1.630000 ;
        RECT 4.445000 1.630000 5.655000 1.780000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.634300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.625000 0.635000 1.885000 1.090000 ;
        RECT 1.625000 1.090000 3.655000 1.260000 ;
        RECT 2.265000 1.850000 4.195000 1.950000 ;
        RECT 2.265000 1.950000 5.145000 2.150000 ;
        RECT 2.265000 2.150000 2.875000 2.980000 ;
        RECT 2.555000 0.635000 2.880000 1.090000 ;
        RECT 3.285000 1.260000 3.655000 1.850000 ;
        RECT 4.815000 2.150000 5.145000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.135000  0.350000 0.385000 0.960000 ;
      RECT 0.135000  0.960000 1.455000 1.130000 ;
      RECT 0.435000  1.950000 1.060000 3.245000 ;
      RECT 0.565000  0.085000 0.895000 0.790000 ;
      RECT 1.195000  0.255000 3.380000 0.425000 ;
      RECT 1.195000  0.425000 1.455000 0.790000 ;
      RECT 1.230000  1.950000 1.560000 2.700000 ;
      RECT 1.285000  1.130000 1.455000 1.430000 ;
      RECT 1.285000  1.430000 3.075000 1.680000 ;
      RECT 1.285000  1.680000 1.455000 1.950000 ;
      RECT 1.765000  1.850000 2.095000 3.245000 ;
      RECT 2.055000  0.425000 2.385000 0.920000 ;
      RECT 3.045000  2.320000 4.645000 3.245000 ;
      RECT 3.050000  0.425000 3.380000 0.750000 ;
      RECT 3.050000  0.750000 4.310000 0.920000 ;
      RECT 3.550000  0.085000 3.880000 0.580000 ;
      RECT 3.980000  0.920000 4.310000 0.960000 ;
      RECT 3.980000  0.960000 5.645000 1.130000 ;
      RECT 4.050000  0.330000 4.310000 0.750000 ;
      RECT 4.480000  0.085000 5.145000 0.790000 ;
      RECT 5.315000  0.350000 5.645000 0.960000 ;
      RECT 5.315000  1.950000 5.600000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_hs__nand2b_4
END LIBRARY
