# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__a311o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.450000 7.075000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.245000 1.450000 7.575000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.420000 5.295000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.470000 1.865000 1.800000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.495000 1.470000 0.825000 1.800000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    ANTENNAPARTIALMETALSIDEAREA  1.869000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.095000 0.810000 0.385000 0.855000 ;
        RECT 0.095000 0.855000 2.785000 0.995000 ;
        RECT 0.095000 0.995000 0.385000 1.040000 ;
        RECT 2.495000 0.810000 2.785000 0.855000 ;
        RECT 2.495000 0.995000 2.785000 1.040000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.125000  0.810000 0.355000 1.040000 ;
      RECT 0.125000  1.040000 0.295000 2.360000 ;
      RECT 0.125000  2.360000 1.505000 2.530000 ;
      RECT 0.305000  2.700000 1.535000 2.905000 ;
      RECT 0.305000  2.905000 2.435000 2.980000 ;
      RECT 0.395000  0.085000 0.725000 0.640000 ;
      RECT 0.755000  2.020000 1.165000 2.190000 ;
      RECT 0.905000  0.390000 1.085000 1.130000 ;
      RECT 0.905000  1.130000 2.325000 1.300000 ;
      RECT 0.995000  1.300000 1.165000 2.020000 ;
      RECT 1.205000  2.980000 2.435000 3.075000 ;
      RECT 1.255000  0.085000 1.585000 0.960000 ;
      RECT 1.335000  1.970000 4.305000 2.140000 ;
      RECT 1.335000  2.140000 1.505000 2.360000 ;
      RECT 1.735000  2.310000 1.905000 2.320000 ;
      RECT 1.735000  2.320000 6.090000 2.460000 ;
      RECT 1.735000  2.460000 5.270000 2.490000 ;
      RECT 1.735000  2.490000 1.905000 2.735000 ;
      RECT 1.755000  0.390000 1.935000 1.130000 ;
      RECT 2.055000  1.300000 2.325000 1.320000 ;
      RECT 2.055000  1.320000 3.905000 1.480000 ;
      RECT 2.055000  1.480000 4.645000 1.650000 ;
      RECT 2.105000  2.660000 2.435000 2.905000 ;
      RECT 2.115000  0.085000 2.365000 0.960000 ;
      RECT 2.525000  1.820000 4.305000 1.970000 ;
      RECT 2.525000  2.140000 4.305000 2.150000 ;
      RECT 2.535000  0.390000 2.920000 0.980000 ;
      RECT 2.535000  0.980000 3.745000 1.150000 ;
      RECT 2.625000  2.660000 2.955000 3.245000 ;
      RECT 3.100000  0.085000 3.315000 0.810000 ;
      RECT 3.495000  0.405000 3.745000 0.980000 ;
      RECT 3.525000  2.660000 3.855000 3.245000 ;
      RECT 3.925000  0.085000 4.175000 0.935000 ;
      RECT 3.925000  0.935000 5.175000 1.150000 ;
      RECT 4.175000  1.150000 5.175000 1.185000 ;
      RECT 4.415000  0.505000 4.745000 0.595000 ;
      RECT 4.415000  0.595000 7.105000 0.765000 ;
      RECT 4.425000  2.660000 4.755000 3.245000 ;
      RECT 4.475000  1.650000 4.645000 1.950000 ;
      RECT 4.475000  1.950000 5.715000 2.120000 ;
      RECT 4.940000  2.290000 6.090000 2.320000 ;
      RECT 4.940000  2.490000 5.270000 2.980000 ;
      RECT 5.365000  0.255000 7.535000 0.425000 ;
      RECT 5.470000  2.630000 5.720000 3.245000 ;
      RECT 5.545000  0.935000 6.105000 1.265000 ;
      RECT 5.545000  1.265000 5.715000 1.950000 ;
      RECT 5.920000  1.950000 7.020000 2.120000 ;
      RECT 5.920000  2.120000 6.090000 2.290000 ;
      RECT 5.920000  2.460000 6.090000 2.980000 ;
      RECT 6.285000  0.985000 7.535000 1.245000 ;
      RECT 6.290000  2.290000 6.650000 3.245000 ;
      RECT 6.775000  0.765000 7.105000 0.815000 ;
      RECT 6.850000  2.120000 7.020000 2.980000 ;
      RECT 7.220000  1.950000 7.550000 3.245000 ;
      RECT 7.285000  0.425000 7.535000 0.985000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  0.840000 0.325000 1.010000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  0.840000 2.725000 1.010000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_hs__a311o_4
END LIBRARY
