# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_hs__sdfsbp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.790000 1.585000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.955000 0.350000 14.290000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.535700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.125000 0.350000 12.620000 1.130000 ;
        RECT 12.450000 1.130000 12.620000 1.820000 ;
        RECT 12.450000 1.820000 12.705000 2.980000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.140000 2.765000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 1.450000 2.045000 1.620000 ;
        RECT 0.505000 1.620000 0.835000 1.850000 ;
        RECT 1.795000 1.260000 2.045000 1.450000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAPARTIALMETALSIDEAREA  1.869000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.295000 1.550000 7.585000 1.595000 ;
        RECT 7.295000 1.595000 9.985000 1.735000 ;
        RECT 7.295000 1.735000 7.585000 1.780000 ;
        RECT 9.695000 1.550000 9.985000 1.595000 ;
        RECT 9.695000 1.735000 9.985000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.275000 1.180000 3.715000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
    END
  END VPB
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.115000  0.350000  0.445000 0.950000 ;
      RECT  0.115000  0.950000  1.140000 1.280000 ;
      RECT  0.115000  1.280000  0.335000 2.290000 ;
      RECT  0.115000  2.290000  2.045000 2.460000 ;
      RECT  0.115000  2.460000  0.365000 2.980000 ;
      RECT  0.565000  2.630000  0.895000 3.245000 ;
      RECT  0.615000  0.085000  0.945000 0.780000 ;
      RECT  1.435000  2.630000  2.385000 2.800000 ;
      RECT  1.435000  2.800000  1.945000 2.960000 ;
      RECT  1.505000  0.350000  1.835000 0.920000 ;
      RECT  1.505000  0.920000  2.385000 1.090000 ;
      RECT  1.795000  1.830000  2.045000 2.290000 ;
      RECT  2.215000  1.090000  2.385000 2.320000 ;
      RECT  2.215000  2.320000  4.925000 2.380000 ;
      RECT  2.215000  2.380000  3.795000 2.490000 ;
      RECT  2.215000  2.490000  2.385000 2.630000 ;
      RECT  2.325000  0.085000  2.655000 0.750000 ;
      RECT  2.555000  2.660000  2.820000 3.245000 ;
      RECT  2.935000  0.340000  3.200000 1.010000 ;
      RECT  2.935000  1.010000  3.105000 1.820000 ;
      RECT  2.935000  1.820000  4.215000 1.990000 ;
      RECT  2.935000  1.990000  3.455000 2.150000 ;
      RECT  3.380000  0.085000  3.710000 1.010000 ;
      RECT  3.575000  2.660000  3.905000 3.245000 ;
      RECT  3.625000  2.210000  4.925000 2.320000 ;
      RECT  3.880000  0.255000  5.030000 0.425000 ;
      RECT  3.880000  0.425000  4.210000 1.010000 ;
      RECT  3.885000  1.220000  4.215000 1.820000 ;
      RECT  4.105000  2.550000  4.355000 2.905000 ;
      RECT  4.105000  2.905000  5.810000 3.075000 ;
      RECT  4.420000  0.595000  4.690000 0.925000 ;
      RECT  4.420000  0.925000  4.590000 2.210000 ;
      RECT  4.590000  2.380000  4.925000 2.735000 ;
      RECT  4.760000  1.370000  5.030000 2.040000 ;
      RECT  4.860000  0.425000  5.030000 1.370000 ;
      RECT  5.120000  2.370000  5.450000 2.735000 ;
      RECT  5.200000  0.350000  5.450000 1.350000 ;
      RECT  5.200000  1.350000  7.110000 1.520000 ;
      RECT  5.200000  1.520000  5.370000 2.370000 ;
      RECT  5.540000  1.690000  5.810000 2.020000 ;
      RECT  5.640000  2.020000  5.810000 2.085000 ;
      RECT  5.640000  2.085000  6.765000 2.255000 ;
      RECT  5.640000  2.255000  5.810000 2.905000 ;
      RECT  5.815000  0.735000  6.770000 0.905000 ;
      RECT  5.815000  0.905000  6.485000 1.180000 ;
      RECT  6.020000  0.085000  6.370000 0.565000 ;
      RECT  6.050000  1.690000  7.105000 1.915000 ;
      RECT  6.175000  2.425000  6.425000 3.245000 ;
      RECT  6.595000  2.255000  6.765000 2.905000 ;
      RECT  6.595000  2.905000  7.445000 3.075000 ;
      RECT  6.600000  0.350000  6.930000 0.735000 ;
      RECT  6.725000  1.190000  7.110000 1.350000 ;
      RECT  6.935000  1.915000  7.105000 2.735000 ;
      RECT  6.940000  0.905000  8.165000 1.075000 ;
      RECT  6.940000  1.075000  7.110000 1.190000 ;
      RECT  7.275000  1.950000  8.830000 2.120000 ;
      RECT  7.275000  2.120000  7.445000 2.905000 ;
      RECT  7.295000  1.245000  7.625000 1.780000 ;
      RECT  7.500000  0.085000  8.295000 0.735000 ;
      RECT  7.615000  2.295000  7.785000 3.245000 ;
      RECT  7.835000  1.075000  8.165000 1.450000 ;
      RECT  7.985000  2.290000  8.315000 2.350000 ;
      RECT  7.985000  2.350000  9.830000 2.520000 ;
      RECT  7.985000  2.520000  8.315000 2.755000 ;
      RECT  8.530000  2.690000  8.860000 2.905000 ;
      RECT  8.530000  2.905000 10.380000 3.075000 ;
      RECT  8.660000  1.350000  8.990000 1.680000 ;
      RECT  8.660000  1.680000  8.830000 1.950000 ;
      RECT  8.785000  0.350000  9.380000 1.050000 ;
      RECT  9.045000  1.850000  9.380000 1.950000 ;
      RECT  9.045000  1.950000 10.170000 2.095000 ;
      RECT  9.045000  2.095000 11.280000 2.120000 ;
      RECT  9.045000  2.120000  9.380000 2.180000 ;
      RECT  9.210000  1.050000  9.380000 1.850000 ;
      RECT  9.580000  2.290000  9.830000 2.350000 ;
      RECT  9.580000  2.520000  9.830000 2.735000 ;
      RECT  9.620000  0.900000 11.395000 1.070000 ;
      RECT  9.620000  1.070000  9.950000 1.230000 ;
      RECT  9.725000  1.550000 10.915000 1.780000 ;
      RECT 10.000000  2.120000 11.280000 2.265000 ;
      RECT 10.050000  2.520000 10.380000 2.905000 ;
      RECT 10.285000  0.085000 10.895000 0.680000 ;
      RECT 10.580000  2.520000 10.750000 3.245000 ;
      RECT 10.585000  1.255000 10.915000 1.550000 ;
      RECT 10.585000  1.780000 10.915000 1.925000 ;
      RECT 10.950000  2.520000 11.280000 2.980000 ;
      RECT 11.065000  0.350000 11.395000 0.900000 ;
      RECT 11.110000  1.640000 11.895000 1.970000 ;
      RECT 11.110000  1.970000 11.280000 2.095000 ;
      RECT 11.110000  2.265000 11.280000 2.520000 ;
      RECT 11.225000  1.070000 11.395000 1.300000 ;
      RECT 11.225000  1.300000 12.235000 1.470000 ;
      RECT 11.500000  2.180000 12.235000 2.350000 ;
      RECT 11.500000  2.350000 11.750000 2.980000 ;
      RECT 11.625000  0.085000 11.955000 1.130000 ;
      RECT 11.950000  2.520000 12.280000 3.245000 ;
      RECT 12.065000  1.470000 12.235000 2.180000 ;
      RECT 12.840000  0.540000 13.255000 1.130000 ;
      RECT 13.005000  1.130000 13.255000 1.220000 ;
      RECT 13.005000  1.220000 13.785000 1.550000 ;
      RECT 13.005000  1.550000 13.255000 2.875000 ;
      RECT 13.455000  0.085000 13.785000 1.050000 ;
      RECT 13.455000  1.995000 13.785000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.580000  7.525000 1.750000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.580000  9.925000 1.750000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
  END
END sky130_fd_sc_hs__sdfsbp_1
END LIBRARY
